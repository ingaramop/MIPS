`timescale 1ns / 1ps

module addPc(input [9:0]inPc, output [9:0]outPc
    );

assign outPc= inPc+1;

endmodule
